`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/19/2021 04:42:00 PM
// Design Name: 
// Module Name: bram_dram_mover_v1_0_S00_AXI_FROM_PS
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bram_dram_mover_v1_0_S00_AXI_FROM_PS(

    );
endmodule
